// platform.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module platform (
		input  wire [7:0]  button_export,             //         button.export
		input  wire        clk_clk,                   //            clk.clk
		inout  wire [15:0] external_flash_data_cf,    // external_flash.data_cf
		output wire        external_flash_we_n,       //               .we_n
		output wire        external_flash_rfu,        //               .rfu
		output wire        external_flash_reset_n_cf, //               .reset_n_cf
		output wire        external_flash_power,      //               .power
		output wire        external_flash_iowr_n,     //               .iowr_n
		output wire        external_flash_iord_n,     //               .iord_n
		output wire [1:0]  external_flash_cs_n,       //               .cs_n
		output wire [10:0] external_flash_addr,       //               .addr
		input  wire        external_flash_iordy,      //               .iordy
		input  wire        external_flash_intrq,      //               .intrq
		input  wire        external_flash_detect_n,   //               .detect_n
		output wire        external_flash_atasel_n,   //               .atasel_n
		output wire        flash_as_dclk,             //       flash_as.dclk
		output wire        flash_as_sce,              //               .sce
		output wire        flash_as_sdo,              //               .sdo
		input  wire        flash_as_data0,            //               .data0
		output wire [7:0]  led_export,                //            led.export
		output wire [31:0] registerdata_readdata,     //   registerdata.readdata
		input  wire        reset_reset_n              //          reset.reset_n
	);

	wire  [31:0] nios_data_master_readdata;                                              // mm_interconnect_0:nios_data_master_readdata -> nios:d_readdata
	wire         nios_data_master_waitrequest;                                           // mm_interconnect_0:nios_data_master_waitrequest -> nios:d_waitrequest
	wire         nios_data_master_debugaccess;                                           // nios:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_data_master_debugaccess
	wire  [16:0] nios_data_master_address;                                               // nios:d_address -> mm_interconnect_0:nios_data_master_address
	wire   [3:0] nios_data_master_byteenable;                                            // nios:d_byteenable -> mm_interconnect_0:nios_data_master_byteenable
	wire         nios_data_master_read;                                                  // nios:d_read -> mm_interconnect_0:nios_data_master_read
	wire         nios_data_master_readdatavalid;                                         // mm_interconnect_0:nios_data_master_readdatavalid -> nios:d_readdatavalid
	wire         nios_data_master_write;                                                 // nios:d_write -> mm_interconnect_0:nios_data_master_write
	wire  [31:0] nios_data_master_writedata;                                             // nios:d_writedata -> mm_interconnect_0:nios_data_master_writedata
	wire  [31:0] nios_instruction_master_readdata;                                       // mm_interconnect_0:nios_instruction_master_readdata -> nios:i_readdata
	wire         nios_instruction_master_waitrequest;                                    // mm_interconnect_0:nios_instruction_master_waitrequest -> nios:i_waitrequest
	wire  [16:0] nios_instruction_master_address;                                        // nios:i_address -> mm_interconnect_0:nios_instruction_master_address
	wire         nios_instruction_master_read;                                           // nios:i_read -> mm_interconnect_0:nios_instruction_master_read
	wire         nios_instruction_master_readdatavalid;                                  // mm_interconnect_0:nios_instruction_master_readdatavalid -> nios:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                 // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;              // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_register0_avalon_slave_0_chipselect;                  // mm_interconnect_0:register0_avalon_slave_0_chipselect -> register0:chipSelect
	wire  [31:0] mm_interconnect_0_register0_avalon_slave_0_readdata;                    // register0:readdata -> mm_interconnect_0:register0_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_register0_avalon_slave_0_address;                     // mm_interconnect_0:register0_avalon_slave_0_address -> register0:address
	wire         mm_interconnect_0_register0_avalon_slave_0_read;                        // mm_interconnect_0:register0_avalon_slave_0_read -> register0:read
	wire         mm_interconnect_0_register0_avalon_slave_0_write;                       // mm_interconnect_0:register0_avalon_slave_0_write -> register0:write
	wire  [31:0] mm_interconnect_0_register0_avalon_slave_0_writedata;                   // mm_interconnect_0:register0_avalon_slave_0_writedata -> register0:writedata
	wire         mm_interconnect_0_external_flash_ctl_chipselect;                        // mm_interconnect_0:external_flash_ctl_chipselect -> external_flash:av_ctl_chipselect_n
	wire   [3:0] mm_interconnect_0_external_flash_ctl_readdata;                          // external_flash:av_ctl_readdata -> mm_interconnect_0:external_flash_ctl_readdata
	wire   [1:0] mm_interconnect_0_external_flash_ctl_address;                           // mm_interconnect_0:external_flash_ctl_address -> external_flash:av_ctl_address
	wire         mm_interconnect_0_external_flash_ctl_read;                              // mm_interconnect_0:external_flash_ctl_read -> external_flash:av_ctl_read_n
	wire         mm_interconnect_0_external_flash_ctl_write;                             // mm_interconnect_0:external_flash_ctl_write -> external_flash:av_ctl_write_n
	wire   [3:0] mm_interconnect_0_external_flash_ctl_writedata;                         // mm_interconnect_0:external_flash_ctl_writedata -> external_flash:av_ctl_writedata
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_readdata;                        // nios:debug_mem_slave_readdata -> mm_interconnect_0:nios_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_debug_mem_slave_waitrequest;                     // nios:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_debug_mem_slave_debugaccess;                     // mm_interconnect_0:nios_debug_mem_slave_debugaccess -> nios:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_debug_mem_slave_address;                         // mm_interconnect_0:nios_debug_mem_slave_address -> nios:debug_mem_slave_address
	wire         mm_interconnect_0_nios_debug_mem_slave_read;                            // mm_interconnect_0:nios_debug_mem_slave_read -> nios:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_debug_mem_slave_byteenable;                      // mm_interconnect_0:nios_debug_mem_slave_byteenable -> nios:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_debug_mem_slave_write;                           // mm_interconnect_0:nios_debug_mem_slave_write -> nios:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_debug_mem_slave_writedata;                       // mm_interconnect_0:nios_debug_mem_slave_writedata -> nios:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_chipselect -> epcs_flash_controller_0:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata;   // epcs_flash_controller_0:readdata -> mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_address -> epcs_flash_controller_0:address
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_read -> epcs_flash_controller_0:read_n
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_write -> epcs_flash_controller_0:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_writedata -> epcs_flash_controller_0:writedata
	wire         mm_interconnect_0_external_flash_ide_chipselect;                        // mm_interconnect_0:external_flash_ide_chipselect -> external_flash:av_ide_chipselect_n
	wire  [15:0] mm_interconnect_0_external_flash_ide_readdata;                          // external_flash:av_ide_readdata -> mm_interconnect_0:external_flash_ide_readdata
	wire   [3:0] mm_interconnect_0_external_flash_ide_address;                           // mm_interconnect_0:external_flash_ide_address -> external_flash:av_ide_address
	wire         mm_interconnect_0_external_flash_ide_read;                              // mm_interconnect_0:external_flash_ide_read -> external_flash:av_ide_read_n
	wire         mm_interconnect_0_external_flash_ide_write;                             // mm_interconnect_0:external_flash_ide_write -> external_flash:av_ide_write_n
	wire  [15:0] mm_interconnect_0_external_flash_ide_writedata;                         // mm_interconnect_0:external_flash_ide_writedata -> external_flash:av_ide_writedata
	wire         mm_interconnect_0_led_s1_chipselect;                                    // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                      // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                       // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                                         // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                     // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                          // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                            // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_s1_address;                             // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                          // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                               // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                           // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                               // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire  [31:0] mm_interconnect_0_button_s1_readdata;                                   // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                                    // mm_interconnect_0:button_s1_address -> button:address
	wire         irq_mapper_receiver0_irq;                                               // external_flash:av_ctl_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                               // external_flash:av_ide_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                               // jtag_uart:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                               // epcs_flash_controller_0:irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios_irq_irq;                                                           // irq_mapper:sender_irq -> nios:irq
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [button:reset_n, epcs_flash_controller_0:reset_n, external_flash:av_reset_n, irq_mapper:reset, jtag_uart:rst_n, led:reset_n, mm_interconnect_0:nios_reset_reset_bridge_in_reset_reset, nios:reset_n, onchip_memory:reset, register0:rst_n, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [epcs_flash_controller_0:reset_req, nios:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]

	platform_button button (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_button_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_button_s1_readdata), //                    .readdata
		.in_port  (button_export)                         // external_connection.export
	);

	platform_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk        (clk_clk),                                                                //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                                     //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver3_irq),                                               //               irq.irq
		.dclk       (flash_as_dclk),                                                          //          external.export
		.sce        (flash_as_sce),                                                           //                  .export
		.sdo        (flash_as_sdo),                                                           //                  .export
		.data0      (flash_as_data0)                                                          //                  .export
	);

	platform_external_flash external_flash (
		.clk                 (clk_clk),                                          //      clk.clk
		.data_cf             (external_flash_data_cf),                           // external.export
		.we_n                (external_flash_we_n),                              //         .export
		.rfu                 (external_flash_rfu),                               //         .export
		.reset_n_cf          (external_flash_reset_n_cf),                        //         .export
		.power               (external_flash_power),                             //         .export
		.iowr_n              (external_flash_iowr_n),                            //         .export
		.iord_n              (external_flash_iord_n),                            //         .export
		.cs_n                (external_flash_cs_n),                              //         .export
		.addr                (external_flash_addr),                              //         .export
		.iordy               (external_flash_iordy),                             //         .export
		.intrq               (external_flash_intrq),                             //         .export
		.detect_n            (external_flash_detect_n),                          //         .export
		.atasel_n            (external_flash_atasel_n),                          //         .export
		.av_reset_n          (~rst_controller_reset_out_reset),                  //    reset.reset_n
		.av_ide_chipselect_n (~mm_interconnect_0_external_flash_ide_chipselect), //      ide.chipselect_n
		.av_ide_read_n       (~mm_interconnect_0_external_flash_ide_read),       //         .read_n
		.av_ide_write_n      (~mm_interconnect_0_external_flash_ide_write),      //         .write_n
		.av_ide_writedata    (mm_interconnect_0_external_flash_ide_writedata),   //         .writedata
		.av_ide_address      (mm_interconnect_0_external_flash_ide_address),     //         .address
		.av_ide_readdata     (mm_interconnect_0_external_flash_ide_readdata),    //         .readdata
		.av_ide_irq          (irq_mapper_receiver1_irq),                         //  ide_irq.irq
		.av_ctl_irq          (irq_mapper_receiver0_irq),                         //  ctl_irq.irq
		.av_ctl_address      (mm_interconnect_0_external_flash_ctl_address),     //      ctl.address
		.av_ctl_chipselect_n (~mm_interconnect_0_external_flash_ctl_chipselect), //         .chipselect_n
		.av_ctl_read_n       (~mm_interconnect_0_external_flash_ctl_read),       //         .read_n
		.av_ctl_write_n      (~mm_interconnect_0_external_flash_ctl_write),      //         .write_n
		.av_ctl_readdata     (mm_interconnect_0_external_flash_ctl_readdata),    //         .readdata
		.av_ctl_writedata    (mm_interconnect_0_external_flash_ctl_writedata)    //         .writedata
	);

	platform_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                   //               irq.irq
	);

	platform_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	platform_nios nios (
		.clk                                 (clk_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                    //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                 //                          .reset_req
		.d_address                           (nios_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_data_master_read),                              //                          .read
		.d_readdata                          (nios_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_data_master_write),                             //                          .write
		.d_writedata                         (nios_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                   //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                    // custom_instruction_master.readra
	);

	platform_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	apexRegister_avalon_interface register0 (
		.clk        (clk_clk),                                               //          clock.clk
		.read       (mm_interconnect_0_register0_avalon_slave_0_read),       // avalon_slave_0.read
		.write      (mm_interconnect_0_register0_avalon_slave_0_write),      //               .write
		.chipSelect (mm_interconnect_0_register0_avalon_slave_0_chipselect), //               .chipselect
		.address    (mm_interconnect_0_register0_avalon_slave_0_address),    //               .address
		.writedata  (mm_interconnect_0_register0_avalon_slave_0_writedata),  //               .writedata
		.readdata   (mm_interconnect_0_register0_avalon_slave_0_readdata),   //               .readdata
		.rst_n      (~rst_controller_reset_out_reset),                       //     reset_sink.reset_n
		.Q          (registerdata_readdata)                                  //       Q_export.readdata
	);

	platform_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                          (clk_clk),                                                                //                                   clk_clk.clk
		.nios_reset_reset_bridge_in_reset_reset               (rst_controller_reset_out_reset),                                         //          nios_reset_reset_bridge_in_reset.reset
		.nios_data_master_address                             (nios_data_master_address),                                               //                          nios_data_master.address
		.nios_data_master_waitrequest                         (nios_data_master_waitrequest),                                           //                                          .waitrequest
		.nios_data_master_byteenable                          (nios_data_master_byteenable),                                            //                                          .byteenable
		.nios_data_master_read                                (nios_data_master_read),                                                  //                                          .read
		.nios_data_master_readdata                            (nios_data_master_readdata),                                              //                                          .readdata
		.nios_data_master_readdatavalid                       (nios_data_master_readdatavalid),                                         //                                          .readdatavalid
		.nios_data_master_write                               (nios_data_master_write),                                                 //                                          .write
		.nios_data_master_writedata                           (nios_data_master_writedata),                                             //                                          .writedata
		.nios_data_master_debugaccess                         (nios_data_master_debugaccess),                                           //                                          .debugaccess
		.nios_instruction_master_address                      (nios_instruction_master_address),                                        //                   nios_instruction_master.address
		.nios_instruction_master_waitrequest                  (nios_instruction_master_waitrequest),                                    //                                          .waitrequest
		.nios_instruction_master_read                         (nios_instruction_master_read),                                           //                                          .read
		.nios_instruction_master_readdata                     (nios_instruction_master_readdata),                                       //                                          .readdata
		.nios_instruction_master_readdatavalid                (nios_instruction_master_readdatavalid),                                  //                                          .readdatavalid
		.button_s1_address                                    (mm_interconnect_0_button_s1_address),                                    //                                 button_s1.address
		.button_s1_readdata                                   (mm_interconnect_0_button_s1_readdata),                                   //                                          .readdata
		.epcs_flash_controller_0_epcs_control_port_address    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_flash_controller_0_epcs_control_port.address
		.epcs_flash_controller_0_epcs_control_port_write      (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),      //                                          .write
		.epcs_flash_controller_0_epcs_control_port_read       (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),       //                                          .read
		.epcs_flash_controller_0_epcs_control_port_readdata   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                                          .readdata
		.epcs_flash_controller_0_epcs_control_port_writedata  (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                                          .writedata
		.epcs_flash_controller_0_epcs_control_port_chipselect (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                                          .chipselect
		.external_flash_ctl_address                           (mm_interconnect_0_external_flash_ctl_address),                           //                        external_flash_ctl.address
		.external_flash_ctl_write                             (mm_interconnect_0_external_flash_ctl_write),                             //                                          .write
		.external_flash_ctl_read                              (mm_interconnect_0_external_flash_ctl_read),                              //                                          .read
		.external_flash_ctl_readdata                          (mm_interconnect_0_external_flash_ctl_readdata),                          //                                          .readdata
		.external_flash_ctl_writedata                         (mm_interconnect_0_external_flash_ctl_writedata),                         //                                          .writedata
		.external_flash_ctl_chipselect                        (mm_interconnect_0_external_flash_ctl_chipselect),                        //                                          .chipselect
		.external_flash_ide_address                           (mm_interconnect_0_external_flash_ide_address),                           //                        external_flash_ide.address
		.external_flash_ide_write                             (mm_interconnect_0_external_flash_ide_write),                             //                                          .write
		.external_flash_ide_read                              (mm_interconnect_0_external_flash_ide_read),                              //                                          .read
		.external_flash_ide_readdata                          (mm_interconnect_0_external_flash_ide_readdata),                          //                                          .readdata
		.external_flash_ide_writedata                         (mm_interconnect_0_external_flash_ide_writedata),                         //                                          .writedata
		.external_flash_ide_chipselect                        (mm_interconnect_0_external_flash_ide_chipselect),                        //                                          .chipselect
		.jtag_uart_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                  //               jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                    //                                          .write
		.jtag_uart_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                     //                                          .read
		.jtag_uart_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                 //                                          .readdata
		.jtag_uart_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                //                                          .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),              //                                          .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),               //                                          .chipselect
		.led_s1_address                                       (mm_interconnect_0_led_s1_address),                                       //                                    led_s1.address
		.led_s1_write                                         (mm_interconnect_0_led_s1_write),                                         //                                          .write
		.led_s1_readdata                                      (mm_interconnect_0_led_s1_readdata),                                      //                                          .readdata
		.led_s1_writedata                                     (mm_interconnect_0_led_s1_writedata),                                     //                                          .writedata
		.led_s1_chipselect                                    (mm_interconnect_0_led_s1_chipselect),                                    //                                          .chipselect
		.nios_debug_mem_slave_address                         (mm_interconnect_0_nios_debug_mem_slave_address),                         //                      nios_debug_mem_slave.address
		.nios_debug_mem_slave_write                           (mm_interconnect_0_nios_debug_mem_slave_write),                           //                                          .write
		.nios_debug_mem_slave_read                            (mm_interconnect_0_nios_debug_mem_slave_read),                            //                                          .read
		.nios_debug_mem_slave_readdata                        (mm_interconnect_0_nios_debug_mem_slave_readdata),                        //                                          .readdata
		.nios_debug_mem_slave_writedata                       (mm_interconnect_0_nios_debug_mem_slave_writedata),                       //                                          .writedata
		.nios_debug_mem_slave_byteenable                      (mm_interconnect_0_nios_debug_mem_slave_byteenable),                      //                                          .byteenable
		.nios_debug_mem_slave_waitrequest                     (mm_interconnect_0_nios_debug_mem_slave_waitrequest),                     //                                          .waitrequest
		.nios_debug_mem_slave_debugaccess                     (mm_interconnect_0_nios_debug_mem_slave_debugaccess),                     //                                          .debugaccess
		.onchip_memory_s1_address                             (mm_interconnect_0_onchip_memory_s1_address),                             //                          onchip_memory_s1.address
		.onchip_memory_s1_write                               (mm_interconnect_0_onchip_memory_s1_write),                               //                                          .write
		.onchip_memory_s1_readdata                            (mm_interconnect_0_onchip_memory_s1_readdata),                            //                                          .readdata
		.onchip_memory_s1_writedata                           (mm_interconnect_0_onchip_memory_s1_writedata),                           //                                          .writedata
		.onchip_memory_s1_byteenable                          (mm_interconnect_0_onchip_memory_s1_byteenable),                          //                                          .byteenable
		.onchip_memory_s1_chipselect                          (mm_interconnect_0_onchip_memory_s1_chipselect),                          //                                          .chipselect
		.onchip_memory_s1_clken                               (mm_interconnect_0_onchip_memory_s1_clken),                               //                                          .clken
		.register0_avalon_slave_0_address                     (mm_interconnect_0_register0_avalon_slave_0_address),                     //                  register0_avalon_slave_0.address
		.register0_avalon_slave_0_write                       (mm_interconnect_0_register0_avalon_slave_0_write),                       //                                          .write
		.register0_avalon_slave_0_read                        (mm_interconnect_0_register0_avalon_slave_0_read),                        //                                          .read
		.register0_avalon_slave_0_readdata                    (mm_interconnect_0_register0_avalon_slave_0_readdata),                    //                                          .readdata
		.register0_avalon_slave_0_writedata                   (mm_interconnect_0_register0_avalon_slave_0_writedata),                   //                                          .writedata
		.register0_avalon_slave_0_chipselect                  (mm_interconnect_0_register0_avalon_slave_0_chipselect)                   //                                          .chipselect
	);

	platform_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios_irq_irq)                    //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
